magic
tech sky130A
magscale 1 2
timestamp 1737921471
<< locali >>
rect 4738 -828 4930 -500
rect 5890 -828 6082 -530
rect 4598 -834 6204 -828
rect 4598 -1014 5128 -834
rect 5308 -1014 6204 -834
rect 4598 -1020 6204 -1014
rect 5890 -1022 6082 -1020
<< viali >>
rect 5128 -1014 5308 -834
<< metal1 >>
rect 4994 2534 5058 2804
rect 4994 1686 5058 1962
rect 4994 846 5058 1120
rect 4994 -6 5058 276
rect 5122 -834 5314 3382
rect 5506 3262 6000 3454
rect 5808 2574 6000 3262
rect 5506 2382 6000 2574
rect 5610 1672 5674 1678
rect 5610 1602 5674 1608
rect 5808 920 6000 2382
rect 5506 728 6000 920
rect 5808 -186 6000 728
rect 5503 -378 6000 -186
rect 5808 -382 6000 -378
rect 5122 -1014 5128 -834
rect 5308 -1014 5314 -834
rect 5122 -1026 5314 -1014
<< via1 >>
rect 4994 1608 5058 1672
rect 5610 1608 5674 1672
<< metal2 >>
rect 4762 1608 4994 1672
rect 5058 1608 5610 1672
rect 5674 1608 5680 1672
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_ex_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 4834 0 1 -682
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 4834 0 1 2694
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 1 0 4834 0 1 1006
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 4834 0 1 1850
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1734044400
transform 1 0 4834 0 1 162
box -184 -128 1336 928
<< labels >>
flabel metal2 4762 1608 4994 1672 0 FreeSans 1600 0 0 0 IBPS_5U
port 0 nsew
flabel metal1 5808 -382 6000 3454 0 FreeSans 1600 0 0 0 IBNS_20U
port 1 nsew
flabel locali 4598 -1020 5128 -828 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
<< end >>
